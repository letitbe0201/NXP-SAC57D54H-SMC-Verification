`include "uvm_macros.svh"
`include "smc_intf.sv"
`include "smc_message.sv"
`include "smc_period.sv"
`include "smc_commanddet.sv"
`include "smc_edgedet.sv"
`include "period_counter.sv"
//`include "recirc_sign.sv"
`include "smc_sequence.sv"
`include "smc_sequencer.sv"
`include "smc_driver.sv"
`include "smc_monin.sv"
`include "smc_monout.sv"
`include "smc_agent.sv"
`include "smc_env.sv"
`include "smc_test.sv"
