`include "uvm_macros.svh"
`include "smc_intf.sv"
`include "smc_message.sv"
`include "smc_period.sv"
`include "smc_duty.sv"
`include "commanddet.sv"
`include "control_col.sv"
`include "clk_control.sv"
`include "smc_edgedet.sv"
`include "period_start.sv"
`include "control_values.sv"
`include "smc_pinval.sv"
`include "off_det.sv"
`include "low_det.sv"
`include "high_det.sv"
`include "pwm_left.sv"
`include "pwm_right.sv"
`include "pwm_center.sv"
`include "per_d_comparison.sv"
`include "smc_sequence.sv"
`include "smc_sequencer.sv"
`include "smc_driver.sv"
`include "smc_monin.sv"
`include "smc_monout.sv"
`include "smc_agent.sv"
`include "smc_env.sv"
`include "smc_test.sv"
