`include "uvm_macros.svh"
`include "smc_intf.sv"
`include "smc_message.sv"
`include "smc_period.sv"
`include "smc_commanddet.sv"
`include "control_col.sv"
`include "smc_clk.sv"
`include "smc_edgedet.sv"
`include "smc_period_start.sv"
`include "control_values.sv"
`include "smc_pinval.sv"
`include "off_det.sv"
`include "low_det.sv"
`include "smc_sequence.sv"
`include "smc_sequencer.sv"
`include "smc_driver.sv"
`include "smc_monin.sv"
`include "smc_monout.sv"
`include "smc_agent.sv"
`include "smc_env.sv"
`include "smc_test.sv"
