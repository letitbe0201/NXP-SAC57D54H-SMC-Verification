class smc_driver extends uvm_driver #(in_msg);

	`uvm_component_utils(smc_driver)
	virtual smc_intf intf;
	in_msg msg;

	function new(string name="smc_driver", uvm_component par=null);
		super.new(name, par);
	endfunction : new

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		if (!uvm_config_db #(virtual smc_intf)::get(this, "", "intf", intf))
			`uvm_fatal("SMC DRIVER", "Something wrong in intf config.")
	endfunction : build_phase

	function void connect_phase(uvm_phase phase);
		super.connect_phase(phase);
	endfunction : connect_phase

	task run_phase(uvm_phase phase);
		forever begin
			seq_item_port.get_next_item(msg);
			@(posedge intf.QCLK) begin
				if (intf.QRESET) begin
					intf.QSEL	<= 0;
					intf.QWRITE	<= 0;
					intf.QADDR	<= 0;
					intf.QDATAIN	<= 0;
				end
				repeat (5) @(posedge intf.QCLK);
				intf.QSEL	= 1;
				intf.QWRITE	= 1;
				intf.QADDR	= 7'h 00;
				intf.QDATAIN	= msg.mcper;
				@(posedge intf.QCLK);	
				intf.QADDR	= 7'h 02;
				intf.QDATAIN	= msg.mcctl1;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 03;
				intf.QDATAIN	= msg.mcctl0;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 10;
				intf.QDATAIN	= msg.mccc3;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 11;
				intf.QDATAIN	= msg.mccc2;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 12;
				intf.QDATAIN	= msg.mccc1;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 13;
				intf.QDATAIN	= msg.mccc0;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 14;
				intf.QDATAIN	= msg.mccc7;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 15;
				intf.QDATAIN	= msg.mccc6;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 16;
				intf.QDATAIN	= msg.mccc5;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 17;
				intf.QDATAIN	= msg.mccc4;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 18;
				intf.QDATAIN	= msg.mccc11;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 19;
				intf.QDATAIN	= msg.mccc10;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1A;
				intf.QDATAIN	= msg.mccc9;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1B;
				intf.QDATAIN	= msg.mccc8;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 20;
				intf.QDATAIN	= msg.mcdc1;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 22;
				intf.QDATAIN	= msg.mcdc0;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 24;
				intf.QDATAIN	= msg.mcdc3;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 26;
				intf.QDATAIN	= msg.mcdc2;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 28;
				intf.QDATAIN	= msg.mcdc5;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2A;
				intf.QDATAIN	= msg.mcdc4;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2C;
				intf.QDATAIN	= msg.mcdc7;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2E;
				intf.QDATAIN	= msg.mcdc6;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 30;
				intf.QDATAIN	= msg.mcdc9;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 32;
				intf.QDATAIN	= msg.mcdc8;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 34;
				intf.QDATAIN	= msg.mcdc11;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 36;
				intf.QDATAIN	= msg.mcdc10;
				@(posedge intf.QCLK);
				intf.QWRITE	= 0;
				intf.QADDR	= 7'h 00 ;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 02;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 03;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 10;
				intf.QDATAIN	= msg.mccc3;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 11;
				intf.QDATAIN	= msg.mccc2;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 12;
				intf.QDATAIN	= msg.mccc1;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 13;
				intf.QDATAIN	= msg.mccc0;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 14;
				intf.QDATAIN	= msg.mccc7;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 15;
				intf.QDATAIN	= msg.mccc6;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 16;
				intf.QDATAIN	= msg.mccc5;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 17;
				intf.QDATAIN	= msg.mccc4;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 18;
				intf.QDATAIN	= msg.mccc11;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 19;
				intf.QDATAIN	= msg.mccc10;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1A;
				intf.QDATAIN	= msg.mccc9;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1B;
				intf.QDATAIN	= msg.mccc8;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 20;
				intf.QDATAIN	= msg.mcdc1;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 22;
				intf.QDATAIN	= msg.mcdc0;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 24;
				intf.QDATAIN	= msg.mcdc3;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 26;
				intf.QDATAIN	= msg.mcdc2;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 28;
				intf.QDATAIN	= msg.mcdc5;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2A;
				intf.QDATAIN	= msg.mcdc4;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2C;
				intf.QDATAIN	= msg.mcdc7;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2E;
				intf.QDATAIN	= msg.mcdc6;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 30;
				intf.QDATAIN	= msg.mcdc9;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 32;
				intf.QDATAIN	= msg.mcdc8;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 34;
				intf.QDATAIN	= msg.mcdc11;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 36;
				intf.QDATAIN	= msg.mcdc10;
				@(posedge intf.QCLK);
				intf.QWRITE	= 0;
				intf.QADDR	= 7'h 00 ;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 02;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 03;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 10;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 11;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 12;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 13;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 14;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 15;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 16;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 17;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 18;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 19;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1A;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 1B;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 20;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 22;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 24;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 26;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 28;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2A;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2C;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 2E;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 30;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 32;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 34;
				@(posedge intf.QCLK);
				intf.QADDR	= 7'h 36;
				@(posedge intf.QCLK);
				intf.QSEL	= 0;
			
			end
			seq_item_port.item_done();
		end
	endtask : run_phase

endclass : smc_driver
